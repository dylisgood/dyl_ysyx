module ysyx_22050854_fetch(
    input clk,
    input rst,
    output [31:0]inst
);

endmodule 